module cpu_add(

);


endmodule