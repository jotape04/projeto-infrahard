module mux_ulaA(
    input wire [31:0] PC,
    output wire [31:0] Data_out
)