module mux_ulaA(
    input wire selector,
    input wire [31:0] PC,
    input wire [31:0] Reg_A,
    input wire [31:0] MDR,
    output wire [31:0] Scr_A
);

    assign Scr_A = {} 

endmodule